module Mode0(
	input control_word_loaded,
	input[2:0] gate);
// we have 3 independent couters, each of which has a mode of operation:


endmodule;